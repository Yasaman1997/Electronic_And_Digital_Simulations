** Profile: "SCHEMATIC1-test"  [ D:\ORCADPROJECTS\Q6\q6-schematic1-test.sim ] 

** Creating circuit file "q6-schematic1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\q6.lib" 
* From [PSPICE NETLIST] section of D:\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM a 0 2.5 0.05 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q6-SCHEMATIC1.net" 


.END
