** Profile: "SCHEMATIC1-1st run"  [ D:\A\e, sources\Electronic\Homeworks\Midterm Project\mid_project\2\2-schematic1-1st run.sim ] 

** Creating circuit file "2-schematic1-1st run.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 4ms 0 4m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\2-SCHEMATIC1.net" 


.END
