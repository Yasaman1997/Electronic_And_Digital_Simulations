** Profile: "SCHEMATIC1- R-2R DAC"  [ D:\A\e, sources\Electronic\Homeworks\BP_Project\BP_Project\R-2R DAC\r-2r dac-schematic1- r-2r dac.sim ] 

** Creating circuit file "r-2r dac-schematic1- r-2r dac.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10000ns 0 100ns 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\r-2r dac-SCHEMATIC1.net" 


.END
