** Profile: "SCHEMATIC1-2nd run"  [ D:\A\e, sources\Electronic\Homeworks\Midterm Project\mid_project\3\3-schematic1-2nd run.sim ] 

** Creating circuit file "3-schematic1-2nd run.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\3-SCHEMATIC1.net" 


.END
