** Profile: "SCHEMATIC1-BinaryWeighted Resistor Ladder DAC"  [ D:\A\e, sources\Electronic\Homeworks\BP_Project\BP_Project\BinaryWeighted Resistor Ladder DAC\binaryweighted resistor ladder dac-schematic1-binaryweighted resistor ladder dac.sim ] 

** Creating circuit file "binaryweighted resistor ladder dac-schematic1-binaryweighted resistor ladder dac.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\binaryweighted resistor ladder dac-SCHEMATIC1.net" 


.END
