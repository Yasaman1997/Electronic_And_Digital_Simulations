** Profile: "SCHEMATIC1-1"  [ D:\DIGITAL_E\HW3_2\ORCAD_SIMULATION_Q11\Q14\q4-schematic1-1.sim ] 

** Creating circuit file "q4-schematic1-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\q4.lib" 
* From [PSPICE NETLIST] section of D:\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM a 0 2.5 0.0005 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q4-SCHEMATIC1.net" 


.END
