** Profile: "SCHEMATIC1-a"  [ D:\A\e, sources\Electronic\Homeworks\BP_Project\BP_Project\A\part_a-schematic1-a.sim ] 

** Creating circuit file "part_a-schematic1-a.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\part_a-SCHEMATIC1.net" 


.END
