** Profile: "SCHEMATIC1-Q1_1"  [ D:\A\e, sources\Electronic\Homeworks\Final_Project\9431022_Yasaman_Mirmohammad_finalProject\1\q1-schematic1-q1_1.sim ] 

** Creating circuit file "q1-schematic1-q1_1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\q1.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ms 0 10us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q1-SCHEMATIC1.net" 


.END
