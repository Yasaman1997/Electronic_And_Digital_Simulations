** Profile: "SCHEMATIC1-Q2"  [ D:\A\e, sources\Electronic\Homeworks\Final_Project\9431022_Yasaman_Mirmohammad_finalProject\2\q2-schematic1-q2.sim ] 

** Creating circuit file "q2-schematic1-q2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ms 0 10us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q2-SCHEMATIC1.net" 


.END
