** Profile: "SCHEMATIC1-1st_run"  [ D:\A\e, sources\Electronic\Homeworks\Midterm Project\mid_project\4\4_2\4-2-schematic1-1st_run.sim ] 

** Creating circuit file "4-2-schematic1-1st_run.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\4-2-SCHEMATIC1.net" 


.END
