** Profile: "SCHEMATIC1-1st run "  [ D:\A\e, sources\Electronic\Homeworks\Midterm Project\mid_project\1\1-schematic1-1st run .sim ] 

** Creating circuit file "1-schematic1-1st run .sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 10 0.01 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\1-SCHEMATIC1.net" 


.END
