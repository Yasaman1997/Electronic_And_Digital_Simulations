** Profile: "SCHEMATIC1-test"  [ D:\DIGITAL_E\HW3_2\ORCAD_SIMULATION_Q11\Q15\q15-SCHEMATIC1-test.sim ] 

** Creating circuit file "q15-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\q15.lib" 
* From [PSPICE NETLIST] section of D:\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM a 0 2.5 0.01 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q15-SCHEMATIC1.net" 


.END
